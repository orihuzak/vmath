module vmath

fn test_fract() {
	assert fract(3.4) == 0.3999999999999999
}
